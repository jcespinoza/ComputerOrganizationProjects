module adder(
    input [3:0] in_value,
    output [3:0] out_value
    );

	assign out_value = in_value + 2;
endmodule
